package test_pkg;
    `include "transaction.svh"
    `include "generator.svh"
    `include "driver.svh"
    `include "monitor.svh"
    `include "coverage.svh"
    `include "scoreboard.svh"
    `include "environment.svh"
//    `include "testbench.svh"
endpackage : test_pkg